package my_pkg;
 import uvm_pkg::*;
`include "mem_seq_item.svh"
`include "mem_sequence.svh"
`include "mem_sequncer.svh"
`include "mem_driver.svh"
`include "mem_monitor.svh"
`include "mem_agent.svh"
`include "mem_scoreboard.svh"
`include "mem_env.svh"
`include "mem_test.svh"
endpackage